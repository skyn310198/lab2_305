library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;

entity test_counter_2 is
end entity test_counter_2;

architecture test of test_counter_2 is
  signal t_Clk, t_Enable, t_Direction, t_Init : std_logic;
  signal t_Q : std_logic_vector(3 downto 0);
  
  
component BCD_counter is
  port(
       Clk, Enable, Direction, Init : in std_logic;
       Q : out std_logic_vector(3 downto 0));
end component BCD_counter;

begin
 DUT: BCD_counter
      port map(t_Clk,t_Enable,t_Direction,t_Init,t_Q);
      
init: process
begin
 t_Direction <= '0','1' after 100 ns,'0' after 200 ns, '1' after 300 ns;
 t_Enable <= '1';
 t_Init <= '0','1' after 50 ns,'0' after 100 ns;
 wait;
end process init;

clk_gen: process
begin
 wait for 5 ns;
 t_Clk <= '1';
 wait for 5 ns;
 t_Clk <= '0';
end process clk_gen;
end architecture test;
